

module top(
    input wire gpio_2
);
wire clk;



endmodule